magic
tech scmos
timestamp 1597030855
<< nwell >>
rect -22 2 17 26
<< polysilicon >>
rect -12 14 -10 16
rect -4 14 -2 16
rect 4 14 6 16
rect -12 0 -10 7
rect -11 -4 -10 0
rect -12 -22 -10 -4
rect -4 -7 -2 7
rect -3 -11 -2 -7
rect -4 -22 -2 -11
rect 4 -14 6 7
rect 5 -18 6 -14
rect 4 -22 6 -18
rect -12 -28 -10 -26
rect -4 -28 -2 -26
rect 4 -28 6 -26
<< ndiffusion >>
rect -15 -26 -12 -22
rect -10 -26 -4 -22
rect -2 -26 4 -22
rect 6 -26 8 -22
<< pdiffusion >>
rect -13 7 -12 14
rect -10 7 -9 14
rect -5 7 -4 14
rect -2 7 -1 14
rect 3 7 4 14
rect 6 7 8 14
<< metal1 >>
rect -22 23 17 26
rect -22 19 -17 23
rect -13 19 -9 23
rect -5 19 -1 23
rect 3 19 8 23
rect 12 19 17 23
rect -22 17 17 19
rect -17 14 -13 17
rect -1 14 3 17
rect -8 0 -5 7
rect 8 0 12 7
rect -24 -4 -15 0
rect -8 -4 12 0
rect -24 -11 -7 -7
rect -24 -18 1 -14
rect 8 -22 12 -4
rect -19 -29 -15 -26
rect -24 -30 17 -29
rect -24 -34 -19 -30
rect -15 -34 -10 -30
rect -6 -34 -1 -30
rect 3 -34 17 -30
rect -24 -35 17 -34
<< ntransistor >>
rect -12 -26 -10 -22
rect -4 -26 -2 -22
rect 4 -26 6 -22
<< ptransistor >>
rect -12 7 -10 14
rect -4 7 -2 14
rect 4 7 6 14
<< polycontact >>
rect -15 -4 -11 0
rect -7 -11 -3 -7
rect 1 -18 5 -14
<< ndcontact >>
rect -19 -26 -15 -22
rect 8 -26 12 -22
<< pdcontact >>
rect -17 7 -13 14
rect -9 7 -5 14
rect -1 7 3 14
rect 8 7 12 14
<< psubstratepcontact >>
rect -19 -34 -15 -30
rect -10 -34 -6 -30
rect -1 -34 3 -30
<< nsubstratencontact >>
rect -17 19 -13 23
rect -9 19 -5 23
rect -1 19 3 23
rect 8 19 12 23
<< labels >>
rlabel metal1 7 -35 11 -33 1 GND
rlabel metal1 -24 -4 -22 0 3 A
rlabel metal1 -24 -11 -22 -7 3 B
rlabel metal1 -24 -18 -22 -14 3 C
rlabel metal1 8 -11 12 -8 1 OUT
rlabel metal1 8 24 12 26 5 VDD
<< end >>
